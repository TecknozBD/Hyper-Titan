module dummy_rtl;

  initial begin
    $display("This is a dummy RTL file.");
  end

endmodule
