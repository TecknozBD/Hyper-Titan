initial begin
  $display("This is a dummy TB file.");
  #10ns;
  $finish;
end
