package dummy_pkg;

  function automatic void dummy_function();
    $display("This is a dummy package function.");
  endfunction
  
endpackage