module hyper_titan_tb;

  rvvcoreminiaxi u_e_core (
      .io_aclk                               ('0),
      .io_aresetn                            ('0),
      .io_axi_slave_write_addr_ready         (),
      .io_axi_slave_write_addr_valid         ('0),
      .io_axi_slave_write_addr_bits_addr     ('0),
      .io_axi_slave_write_addr_bits_prot     ('0),
      .io_axi_slave_write_addr_bits_id       ('0),
      .io_axi_slave_write_addr_bits_len      ('0),
      .io_axi_slave_write_addr_bits_size     ('0),
      .io_axi_slave_write_addr_bits_burst    ('0),
      .io_axi_slave_write_addr_bits_lock     ('0),
      .io_axi_slave_write_addr_bits_cache    ('0),
      .io_axi_slave_write_addr_bits_qos      ('0),
      .io_axi_slave_write_addr_bits_region   ('0),
      .io_axi_slave_write_data_ready         (),
      .io_axi_slave_write_data_valid         ('0),
      .io_axi_slave_write_data_bits_data     ('0),
      .io_axi_slave_write_data_bits_last     ('0),
      .io_axi_slave_write_data_bits_strb     ('0),
      .io_axi_slave_write_resp_ready         ('0),
      .io_axi_slave_write_resp_valid         (),
      .io_axi_slave_write_resp_bits_id       (),
      .io_axi_slave_write_resp_bits_resp     (),
      .io_axi_slave_read_addr_ready          (),
      .io_axi_slave_read_addr_valid          ('0),
      .io_axi_slave_read_addr_bits_addr      ('0),
      .io_axi_slave_read_addr_bits_prot      ('0),
      .io_axi_slave_read_addr_bits_id        ('0),
      .io_axi_slave_read_addr_bits_len       ('0),
      .io_axi_slave_read_addr_bits_size      ('0),
      .io_axi_slave_read_addr_bits_burst     ('0),
      .io_axi_slave_read_addr_bits_lock      ('0),
      .io_axi_slave_read_addr_bits_cache     ('0),
      .io_axi_slave_read_addr_bits_qos       ('0),
      .io_axi_slave_read_addr_bits_region    ('0),
      .io_axi_slave_read_data_ready          ('0),
      .io_axi_slave_read_data_valid          (),
      .io_axi_slave_read_data_bits_data      (),
      .io_axi_slave_read_data_bits_id        (),
      .io_axi_slave_read_data_bits_resp      (),
      .io_axi_slave_read_data_bits_last      (),
      .io_axi_master_write_addr_ready        ('0),
      .io_axi_master_write_addr_valid        (),
      .io_axi_master_write_addr_bits_addr    (),
      .io_axi_master_write_addr_bits_prot    (),
      .io_axi_master_write_addr_bits_id      (),
      .io_axi_master_write_addr_bits_len     (),
      .io_axi_master_write_addr_bits_size    (),
      .io_axi_master_write_addr_bits_burst   (),
      .io_axi_master_write_addr_bits_lock    (),
      .io_axi_master_write_addr_bits_cache   (),
      .io_axi_master_write_addr_bits_qos     (),
      .io_axi_master_write_addr_bits_region  (),
      .io_axi_master_write_data_ready        ('0),
      .io_axi_master_write_data_valid        (),
      .io_axi_master_write_data_bits_data    (),
      .io_axi_master_write_data_bits_last    (),
      .io_axi_master_write_data_bits_strb    (),
      .io_axi_master_write_resp_ready        (),
      .io_axi_master_write_resp_valid        ('0),
      .io_axi_master_write_resp_bits_id      ('0),
      .io_axi_master_write_resp_bits_resp    ('0),
      .io_axi_master_read_addr_ready         ('0),
      .io_axi_master_read_addr_valid         (),
      .io_axi_master_read_addr_bits_addr     (),
      .io_axi_master_read_addr_bits_prot     (),
      .io_axi_master_read_addr_bits_id       (),
      .io_axi_master_read_addr_bits_len      (),
      .io_axi_master_read_addr_bits_size     (),
      .io_axi_master_read_addr_bits_burst    (),
      .io_axi_master_read_addr_bits_lock     (),
      .io_axi_master_read_addr_bits_cache    (),
      .io_axi_master_read_addr_bits_qos      (),
      .io_axi_master_read_addr_bits_region   (),
      .io_axi_master_read_data_ready         (),
      .io_axi_master_read_data_valid         ('0),
      .io_axi_master_read_data_bits_data     ('0),
      .io_axi_master_read_data_bits_id       ('0),
      .io_axi_master_read_data_bits_resp     ('0),
      .io_axi_master_read_data_bits_last     ('0),
      .io_halted                             (),
      .io_fault                              (),
      .io_wfi                                (),
      .io_irq                                ('0),
      .io_debug_en                           (),
      .io_debug_addr_0                       (),
      .io_debug_addr_1                       (),
      .io_debug_addr_2                       (),
      .io_debug_addr_3                       (),
      .io_debug_inst_0                       (),
      .io_debug_inst_1                       (),
      .io_debug_inst_2                       (),
      .io_debug_inst_3                       (),
      .io_debug_cycles                       (),
      .io_debug_dbus_valid                   (),
      .io_debug_dbus_bits_addr               (),
      .io_debug_dbus_bits_wdata              (),
      .io_debug_dbus_bits_write              (),
      .io_debug_dispatch_0_instFire          (),
      .io_debug_dispatch_0_instAddr          (),
      .io_debug_dispatch_0_instInst          (),
      .io_debug_dispatch_1_instFire          (),
      .io_debug_dispatch_1_instAddr          (),
      .io_debug_dispatch_1_instInst          (),
      .io_debug_dispatch_2_instFire          (),
      .io_debug_dispatch_2_instAddr          (),
      .io_debug_dispatch_2_instInst          (),
      .io_debug_dispatch_3_instFire          (),
      .io_debug_dispatch_3_instAddr          (),
      .io_debug_dispatch_3_instInst          (),
      .io_debug_regfile_writeAddr_0_valid    (),
      .io_debug_regfile_writeAddr_0_bits     (),
      .io_debug_regfile_writeAddr_1_valid    (),
      .io_debug_regfile_writeAddr_1_bits     (),
      .io_debug_regfile_writeAddr_2_valid    (),
      .io_debug_regfile_writeAddr_2_bits     (),
      .io_debug_regfile_writeAddr_3_valid    (),
      .io_debug_regfile_writeAddr_3_bits     (),
      .io_debug_regfile_writeData_0_valid    (),
      .io_debug_regfile_writeData_0_bits_addr(),
      .io_debug_regfile_writeData_0_bits_data(),
      .io_debug_regfile_writeData_1_valid    (),
      .io_debug_regfile_writeData_1_bits_addr(),
      .io_debug_regfile_writeData_1_bits_data(),
      .io_debug_regfile_writeData_2_valid    (),
      .io_debug_regfile_writeData_2_bits_addr(),
      .io_debug_regfile_writeData_2_bits_data(),
      .io_debug_regfile_writeData_3_valid    (),
      .io_debug_regfile_writeData_3_bits_addr(),
      .io_debug_regfile_writeData_3_bits_data(),
      .io_debug_regfile_writeData_4_valid    (),
      .io_debug_regfile_writeData_4_bits_addr(),
      .io_debug_regfile_writeData_4_bits_data(),
      .io_debug_regfile_writeData_5_valid    (),
      .io_debug_regfile_writeData_5_bits_addr(),
      .io_debug_regfile_writeData_5_bits_data(),
      .io_debug_float_writeAddr_valid        (),
      .io_debug_float_writeAddr_bits         (),
      .io_debug_float_writeData_0_valid      (),
      .io_debug_float_writeData_0_bits_addr  (),
      .io_debug_float_writeData_0_bits_data  (),
      .io_debug_float_writeData_1_valid      (),
      .io_debug_float_writeData_1_bits_addr  (),
      .io_debug_float_writeData_1_bits_data  (),
      .io_slog_valid                         (),
      .io_slog_addr                          (),
      .io_slog_data                          (),
      .io_te                                 ('0)
  );

  ariane u_p_core (
      .clk_i      ('0),
      .rst_ni     ('0),
      .boot_addr_i('0),
      .hart_id_i  ('0),
      .irq_i      ('0),
      .ipi_i      ('0),
      .time_irq_i ('0),
      .debug_req_i('0),
      .axi_req_o  (),
      .axi_resp_i ('0)
  );

  initial begin
    $display("Test running...");
    #10ns;
    $finish;
  end

endmodule
