interface dummy_if;

  initial begin
    $display("This is a dummy interface.");
  end

endinterface
